library verilog;
use verilog.vl_types.all;
entity AluFinal_vlg_vec_tst is
end AluFinal_vlg_vec_tst;
